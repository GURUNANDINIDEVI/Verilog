module or_gate(
    input wire A,    // Input A
    input wire B,    // Input B
    output wire Y    // Output Y
);

assign Y = A | B;  // OR operation

endmodule
