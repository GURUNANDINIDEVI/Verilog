//T.Guru Nandini Devi
//nandinidevitekumudigmail.com
module binary_multiplier_2bit (
    input  [1:0] A,
    input  [1:0] B,
    output [3:0] Product
);
    assign Product = A * B;
endmodule
