//T.Guru Nandini Devi
//nandinidevitekumudi@gmail.com
module or_gate(
    input wire a,    // Input A
    input wire b,    // Input B
    output wire y    // Output Y
);

assign y = a | b;  // OR operation

endmodule
