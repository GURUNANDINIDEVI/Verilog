//T.Guru Nandini Devi
//nandinidevitekumudi@gmail.com
module clock_buffer (
    input wire clk_in,
    output wire clk_out
);

assign clk_out = clk_in;

endmodule
