//T.Guru Nandini Devi
//nandinidevitekumudi@gmail.com
module square_generator (
    input  [1:0] a,
    output [3:0] square
);

assign square = a * a;

endmodule
