//T.Guru Nandini Devi
//nandinidevitekumudi@gmail.com
module and_gate(
    input wire A,    // Input A
    input wire B,    // Input B
    output wire Y    // Output Y
);

assign Y = A & B;  // AND operation

endmodule
